`ifndef FULL_ADD_V
`define FULL_ADD_V
module full_add(
  input [31:0] a,
  input [31:0] b,
  input c_in,
  output [31:0] sum,
  output c_out
);
wire p0,g0,c0;
wire p1,g1,c1;
wire p2,g2,c2;
wire p3,g3,c3;
wire p4,g4,c4;
wire p5,g5,c5;
wire p6,g6,c6;
wire p7,g7,c7;
wire p8,g8,c8;
wire p9,g9,c9;
wire p10,g10,c10;
wire p11,g11,c11;
wire p12,g12,c12;
wire p13,g13,c13;
wire p14,g14,c14;
wire p15,g15,c15;
wire p16,g16,c16;
wire p17,g17,c17;
wire p18,g18,c18;
wire p19,g19,c19;
wire p20,g20,c20;
wire p21,g21,c21;
wire p22,g22,c22;
wire p23,g23,c23;
wire p24,g24,c24;
wire p25,g25,c25;
wire p26,g26,c26;
wire p27,g27,c27;
wire p28,g28,c28;
wire p29,g29,c29;
wire p30,g30,c30;
wire p31,g31,c31;
wire c32;
assign p0 = a[0] ^ b[0];
assign p1 = a[1] ^ b[1];
assign p2 = a[2] ^ b[2];
assign p3 = a[3] ^ b[3];
assign p4 = a[4] ^ b[4];
assign p5 = a[5] ^ b[5];
assign p6 = a[6] ^ b[6];
assign p7 = a[7] ^ b[7];
assign p8 = a[8] ^ b[8];
assign p9 = a[9] ^ b[9];
assign p10 = a[10] ^ b[10];
assign p11 = a[11] ^ b[11];
assign p12 = a[12] ^ b[12];
assign p13 = a[13] ^ b[13];
assign p14 = a[14] ^ b[14];
assign p15 = a[15] ^ b[15];
assign p16 = a[16] ^ b[16];
assign p17 = a[17] ^ b[17];
assign p18 = a[18] ^ b[18];
assign p19 = a[19] ^ b[19];
assign p20 = a[20] ^ b[20];
assign p21 = a[21] ^ b[21];
assign p22 = a[22] ^ b[22];
assign p23 = a[23] ^ b[23];
assign p24 = a[24] ^ b[24];
assign p25 = a[25] ^ b[25];
assign p26 = a[26] ^ b[26];
assign p27 = a[27] ^ b[27];
assign p28 = a[28] ^ b[28];
assign p29 = a[29] ^ b[29];
assign p30 = a[30] ^ b[30];
assign p31 = a[31] ^ b[31];
assign g0 = a[0] & b[0];
assign g1 = a[1] & b[1];
assign g2 = a[2] & b[2];
assign g3 = a[3] & b[3];
assign g4 = a[4] & b[4];
assign g5 = a[5] & b[5];
assign g6 = a[6] & b[6];
assign g7 = a[7] & b[7];
assign g8 = a[8] & b[8];
assign g9 = a[9] & b[9];
assign g10 = a[10] & b[10];
assign g11 = a[11] & b[11];
assign g12 = a[12] & b[12];
assign g13 = a[13] & b[13];
assign g14 = a[14] & b[14];
assign g15 = a[15] & b[15];
assign g16 = a[16] & b[16];
assign g17 = a[17] & b[17];
assign g18 = a[18] & b[18];
assign g19 = a[19] & b[19];
assign g20 = a[20] & b[20];
assign g21 = a[21] & b[21];
assign g22 = a[22] & b[22];
assign g23 = a[23] & b[23];
assign g24 = a[24] & b[24];
assign g25 = a[25] & b[25];
assign g26 = a[26] & b[26];
assign g27 = a[27] & b[27];
assign g28 = a[28] & b[28];
assign g29 = a[29] & b[29];
assign g30 = a[30] & b[30];
assign g31 = a[31] & b[31];
assign c0 = c_in;
assign c1 = (g0) | (c0 & p0);
assign c2 = (g1) | (g0 & p1) | (c0 & p0 & p1);
assign c3 = (g2) | (g1 & p2) | (g0 & p1 & p2) | (c0 & p0 & p1 & p2);
assign c4 = (g3) | (g2 & p3) | (g1 & p2 & p3) | (g0 & p1 & p2 & p3) | (c0 & p0 & p1 & p2 & p3);
assign c5 = (g4) | (g3 & p4) | (g2 & p3 & p4) | (g1 & p2 & p3 & p4) | (g0 & p1 & p2 & p3 & p4) | (c0 & p0 & p1 & p2 & p3 & p4);
assign c6 = (g5) | (g4 & p5) | (g3 & p4 & p5) | (g2 & p3 & p4 & p5) | (g1 & p2 & p3 & p4 & p5) | (g0 & p1 & p2 & p3 & p4 & p5) | (c0 & p0 & p1 & p2 & p3 & p4 & p5);
assign c7 = (g6) | (g5 & p6) | (g4 & p5 & p6) | (g3 & p4 & p5 & p6) | (g2 & p3 & p4 & p5 & p6) | (g1 & p2 & p3 & p4 & p5 & p6) | (g0 & p1 & p2 & p3 & p4 & p5 & p6) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6);
assign c8 = (g7) | (g6 & p7) | (g5 & p6 & p7) | (g4 & p5 & p6 & p7) | (g3 & p4 & p5 & p6 & p7) | (g2 & p3 & p4 & p5 & p6 & p7) | (g1 & p2 & p3 & p4 & p5 & p6 & p7) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7);
assign c9 = (g8) | (g7 & p8) | (g6 & p7 & p8) | (g5 & p6 & p7 & p8) | (g4 & p5 & p6 & p7 & p8) | (g3 & p4 & p5 & p6 & p7 & p8) | (g2 & p3 & p4 & p5 & p6 & p7 & p8) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8);
assign c10 = (g9) | (g8 & p9) | (g7 & p8 & p9) | (g6 & p7 & p8 & p9) | (g5 & p6 & p7 & p8 & p9) | (g4 & p5 & p6 & p7 & p8 & p9) | (g3 & p4 & p5 & p6 & p7 & p8 & p9) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9);
assign c11 = (g10) | (g9 & p10) | (g8 & p9 & p10) | (g7 & p8 & p9 & p10) | (g6 & p7 & p8 & p9 & p10) | (g5 & p6 & p7 & p8 & p9 & p10) | (g4 & p5 & p6 & p7 & p8 & p9 & p10) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10);
assign c12 = (g11) | (g10 & p11) | (g9 & p10 & p11) | (g8 & p9 & p10 & p11) | (g7 & p8 & p9 & p10 & p11) | (g6 & p7 & p8 & p9 & p10 & p11) | (g5 & p6 & p7 & p8 & p9 & p10 & p11) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11);
assign c13 = (g12) | (g11 & p12) | (g10 & p11 & p12) | (g9 & p10 & p11 & p12) | (g8 & p9 & p10 & p11 & p12) | (g7 & p8 & p9 & p10 & p11 & p12) | (g6 & p7 & p8 & p9 & p10 & p11 & p12) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12);
assign c14 = (g13) | (g12 & p13) | (g11 & p12 & p13) | (g10 & p11 & p12 & p13) | (g9 & p10 & p11 & p12 & p13) | (g8 & p9 & p10 & p11 & p12 & p13) | (g7 & p8 & p9 & p10 & p11 & p12 & p13) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13);
assign c15 = (g14) | (g13 & p14) | (g12 & p13 & p14) | (g11 & p12 & p13 & p14) | (g10 & p11 & p12 & p13 & p14) | (g9 & p10 & p11 & p12 & p13 & p14) | (g8 & p9 & p10 & p11 & p12 & p13 & p14) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14);
assign c16 = (g15) | (g14 & p15) | (g13 & p14 & p15) | (g12 & p13 & p14 & p15) | (g11 & p12 & p13 & p14 & p15) | (g10 & p11 & p12 & p13 & p14 & p15) | (g9 & p10 & p11 & p12 & p13 & p14 & p15) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15);
assign c17 = (g16) | (g15 & p16) | (g14 & p15 & p16) | (g13 & p14 & p15 & p16) | (g12 & p13 & p14 & p15 & p16) | (g11 & p12 & p13 & p14 & p15 & p16) | (g10 & p11 & p12 & p13 & p14 & p15 & p16) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16);
assign c18 = (g17) | (g16 & p17) | (g15 & p16 & p17) | (g14 & p15 & p16 & p17) | (g13 & p14 & p15 & p16 & p17) | (g12 & p13 & p14 & p15 & p16 & p17) | (g11 & p12 & p13 & p14 & p15 & p16 & p17) | (g10 & p11 & p12 & p13 & p14 & p15 & p16 & p17) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17);
assign c19 = (g18) | (g17 & p18) | (g16 & p17 & p18) | (g15 & p16 & p17 & p18) | (g14 & p15 & p16 & p17 & p18) | (g13 & p14 & p15 & p16 & p17 & p18) | (g12 & p13 & p14 & p15 & p16 & p17 & p18) | (g11 & p12 & p13 & p14 & p15 & p16 & p17 & p18) | (g10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18);
assign c20 = (g19) | (g18 & p19) | (g17 & p18 & p19) | (g16 & p17 & p18 & p19) | (g15 & p16 & p17 & p18 & p19) | (g14 & p15 & p16 & p17 & p18 & p19) | (g13 & p14 & p15 & p16 & p17 & p18 & p19) | (g12 & p13 & p14 & p15 & p16 & p17 & p18 & p19) | (g11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19) | (g10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19);
assign c21 = (g20) | (g19 & p20) | (g18 & p19 & p20) | (g17 & p18 & p19 & p20) | (g16 & p17 & p18 & p19 & p20) | (g15 & p16 & p17 & p18 & p19 & p20) | (g14 & p15 & p16 & p17 & p18 & p19 & p20) | (g13 & p14 & p15 & p16 & p17 & p18 & p19 & p20) | (g12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20) | (g11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20) | (g10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20);
assign c22 = (g21) | (g20 & p21) | (g19 & p20 & p21) | (g18 & p19 & p20 & p21) | (g17 & p18 & p19 & p20 & p21) | (g16 & p17 & p18 & p19 & p20 & p21) | (g15 & p16 & p17 & p18 & p19 & p20 & p21) | (g14 & p15 & p16 & p17 & p18 & p19 & p20 & p21) | (g13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21) | (g12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21) | (g11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21) | (g10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21);
assign c23 = (g22) | (g21 & p22) | (g20 & p21 & p22) | (g19 & p20 & p21 & p22) | (g18 & p19 & p20 & p21 & p22) | (g17 & p18 & p19 & p20 & p21 & p22) | (g16 & p17 & p18 & p19 & p20 & p21 & p22) | (g15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (g14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (g13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (g12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (g11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (g10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22);
assign c24 = (g23) | (g22 & p23) | (g21 & p22 & p23) | (g20 & p21 & p22 & p23) | (g19 & p20 & p21 & p22 & p23) | (g18 & p19 & p20 & p21 & p22 & p23) | (g17 & p18 & p19 & p20 & p21 & p22 & p23) | (g16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23);
assign c25 = (g24) | (g23 & p24) | (g22 & p23 & p24) | (g21 & p22 & p23 & p24) | (g20 & p21 & p22 & p23 & p24) | (g19 & p20 & p21 & p22 & p23 & p24) | (g18 & p19 & p20 & p21 & p22 & p23 & p24) | (g17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24);
assign c26 = (g25) | (g24 & p25) | (g23 & p24 & p25) | (g22 & p23 & p24 & p25) | (g21 & p22 & p23 & p24 & p25) | (g20 & p21 & p22 & p23 & p24 & p25) | (g19 & p20 & p21 & p22 & p23 & p24 & p25) | (g18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25);
assign c27 = (g26) | (g25 & p26) | (g24 & p25 & p26) | (g23 & p24 & p25 & p26) | (g22 & p23 & p24 & p25 & p26) | (g21 & p22 & p23 & p24 & p25 & p26) | (g20 & p21 & p22 & p23 & p24 & p25 & p26) | (g19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26);
assign c28 = (g27) | (g26 & p27) | (g25 & p26 & p27) | (g24 & p25 & p26 & p27) | (g23 & p24 & p25 & p26 & p27) | (g22 & p23 & p24 & p25 & p26 & p27) | (g21 & p22 & p23 & p24 & p25 & p26 & p27) | (g20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27);
assign c29 = (g28) | (g27 & p28) | (g26 & p27 & p28) | (g25 & p26 & p27 & p28) | (g24 & p25 & p26 & p27 & p28) | (g23 & p24 & p25 & p26 & p27 & p28) | (g22 & p23 & p24 & p25 & p26 & p27 & p28) | (g21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28);
assign c30 = (g29) | (g28 & p29) | (g27 & p28 & p29) | (g26 & p27 & p28 & p29) | (g25 & p26 & p27 & p28 & p29) | (g24 & p25 & p26 & p27 & p28 & p29) | (g23 & p24 & p25 & p26 & p27 & p28 & p29) | (g22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29);
assign c31 = (g30) | (g29 & p30) | (g28 & p29 & p30) | (g27 & p28 & p29 & p30) | (g26 & p27 & p28 & p29 & p30) | (g25 & p26 & p27 & p28 & p29 & p30) | (g24 & p25 & p26 & p27 & p28 & p29 & p30) | (g23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30);
assign c32 = (g31) | (g30 & p31) | (g29 & p30 & p31) | (g28 & p29 & p30 & p31) | (g27 & p28 & p29 & p30 & p31) | (g26 & p27 & p28 & p29 & p30 & p31) | (g25 & p26 & p27 & p28 & p29 & p30 & p31) | (g24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (g0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31) | (c0 & p0 & p1 & p2 & p3 & p4 & p5 & p6 & p7 & p8 & p9 & p10 & p11 & p12 & p13 & p14 & p15 & p16 & p17 & p18 & p19 & p20 & p21 & p22 & p23 & p24 & p25 & p26 & p27 & p28 & p29 & p30 & p31);
assign sum[0] = p0 ^ c0;
assign sum[1] = p1 ^ c1;
assign sum[2] = p2 ^ c2;
assign sum[3] = p3 ^ c3;
assign sum[4] = p4 ^ c4;
assign sum[5] = p5 ^ c5;
assign sum[6] = p6 ^ c6;
assign sum[7] = p7 ^ c7;
assign sum[8] = p8 ^ c8;
assign sum[9] = p9 ^ c9;
assign sum[10] = p10 ^ c10;
assign sum[11] = p11 ^ c11;
assign sum[12] = p12 ^ c12;
assign sum[13] = p13 ^ c13;
assign sum[14] = p14 ^ c14;
assign sum[15] = p15 ^ c15;
assign sum[16] = p16 ^ c16;
assign sum[17] = p17 ^ c17;
assign sum[18] = p18 ^ c18;
assign sum[19] = p19 ^ c19;
assign sum[20] = p20 ^ c20;
assign sum[21] = p21 ^ c21;
assign sum[22] = p22 ^ c22;
assign sum[23] = p23 ^ c23;
assign sum[24] = p24 ^ c24;
assign sum[25] = p25 ^ c25;
assign sum[26] = p26 ^ c26;
assign sum[27] = p27 ^ c27;
assign sum[28] = p28 ^ c28;
assign sum[29] = p29 ^ c29;
assign sum[30] = p30 ^ c30;
assign sum[31] = p31 ^ c31;
assign c_out = c32;
endmodule
`endif
