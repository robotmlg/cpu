`ifndef MUL_V
`define MUL_V
module mul(
  input [31:0] a,
  input [31:0] b,
  output [63:0] prod
);
wire [63:0] P;
wire [31:0] p0;
wire [31:0] p1;
wire [31:0] p2;
wire [31:0] p3;
wire [31:0] p4;
wire [31:0] p5;
wire [31:0] p6;
wire [31:0] p7;
wire [31:0] p8;
wire [31:0] p9;
wire [31:0] p10;
wire [31:0] p11;
wire [31:0] p12;
wire [31:0] p13;
wire [31:0] p14;
wire [31:0] p15;
wire [31:0] p16;
wire [31:0] p17;
wire [31:0] p18;
wire [31:0] p19;
wire [31:0] p20;
wire [31:0] p21;
wire [31:0] p22;
wire [31:0] p23;
wire [31:0] p24;
wire [31:0] p25;
wire [31:0] p26;
wire [31:0] p27;
wire [31:0] p28;
wire [31:0] p29;
wire [31:0] p30;
wire [31:0] p31;
assign p0 = {32{a[0]}} & b;
assign p1 = {32{a[1]}} & b;
assign p2 = {32{a[2]}} & b;
assign p3 = {32{a[3]}} & b;
assign p4 = {32{a[4]}} & b;
assign p5 = {32{a[5]}} & b;
assign p6 = {32{a[6]}} & b;
assign p7 = {32{a[7]}} & b;
assign p8 = {32{a[8]}} & b;
assign p9 = {32{a[9]}} & b;
assign p10 = {32{a[10]}} & b;
assign p11 = {32{a[11]}} & b;
assign p12 = {32{a[12]}} & b;
assign p13 = {32{a[13]}} & b;
assign p14 = {32{a[14]}} & b;
assign p15 = {32{a[15]}} & b;
assign p16 = {32{a[16]}} & b;
assign p17 = {32{a[17]}} & b;
assign p18 = {32{a[18]}} & b;
assign p19 = {32{a[19]}} & b;
assign p20 = {32{a[20]}} & b;
assign p21 = {32{a[21]}} & b;
assign p22 = {32{a[22]}} & b;
assign p23 = {32{a[23]}} & b;
assign p24 = {32{a[24]}} & b;
assign p25 = {32{a[25]}} & b;
assign p26 = {32{a[26]}} & b;
assign p27 = {32{a[27]}} & b;
assign p28 = {32{a[28]}} & b;
assign p29 = {32{a[29]}} & b;
assign p30 = {32{a[30]}} & b;
assign p31 = {32{a[31]}} & b;
assign P = {1'b1,~p0[31],p0[30:0]} + {~p1[31],p1[30:0],1'b0} + {~p2[31],p2[30:0],2'b0} + {~p3[31],p3[30:0],3'b0} + {~p4[31],p4[30:0],4'b0} + {~p5[31],p5[30:0],5'b0} + {~p6[31],p6[30:0],6'b0} + {~p7[31],p7[30:0],7'b0} + {~p8[31],p8[30:0],8'b0} + {~p9[31],p9[30:0],9'b0} + {~p10[31],p10[30:0],10'b0} + {~p11[31],p11[30:0],11'b0} + {~p12[31],p12[30:0],12'b0} + {~p13[31],p13[30:0],13'b0} + {~p14[31],p14[30:0],14'b0} + {~p15[31],p15[30:0],15'b0} + {~p16[31],p16[30:0],16'b0} + {~p17[31],p17[30:0],17'b0} + {~p18[31],p18[30:0],18'b0} + {~p19[31],p19[30:0],19'b0} + {~p20[31],p20[30:0],20'b0} + {~p21[31],p21[30:0],21'b0} + {~p22[31],p22[30:0],22'b0} + {~p23[31],p23[30:0],23'b0} + {~p24[31],p24[30:0],24'b0} + {~p25[31],p25[30:0],25'b0} + {~p26[31],p26[30:0],26'b0} + {~p27[31],p27[30:0],27'b0} + {~p28[31],p28[30:0],28'b0} + {~p29[31],p29[30:0],29'b0} + {~p30[31],p30[30:0],30'b0} + {1'b1,~p31[31],p31[30],p31[29],p31[28],p31[27],p31[26],p31[25],p31[24],p31[23],p31[22],p31[21],p31[20],p31[19],p31[18],p31[17],p31[16],p31[15],p31[14],p31[13],p31[12],p31[11],p31[10],p31[9],p31[8],p31[7],p31[6],p31[5],p31[4],p31[3],p31[2],p31[1],p31[0],31'b0};
assign prod = P;
endmodule
`endif
